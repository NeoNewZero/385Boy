// nios_system.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module nios_system (
		output wire [15:0] address_export,       //        address.export
		input  wire [3:0]  buttons_export,       //        buttons.export
		input  wire        clk_clk,              //            clk.clk
		input  wire [7:0]  din_export,           //            din.export
		input  wire        gameboy_clk_clk,      //    gameboy_clk.clk
		output wire [7:0]  leds_export,          //           leds.export
		input  wire        reset_reset_n,        //          reset.reset_n
		output wire        sdram_clk_clk,        //      sdram_clk.clk
		output wire [12:0] sdram_wire_addr,      //     sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,        //               .ba
		output wire        sdram_wire_cas_n,     //               .cas_n
		output wire        sdram_wire_cke,       //               .cke
		output wire        sdram_wire_cs_n,      //               .cs_n
		inout  wire [31:0] sdram_wire_dq,        //               .dq
		output wire [3:0]  sdram_wire_dqm,       //               .dqm
		output wire        sdram_wire_ras_n,     //               .ras_n
		output wire        sdram_wire_we_n,      //               .we_n
		inout  wire [15:0] sram_DQ,              //           sram.DQ
		output wire [19:0] sram_ADDR,            //               .ADDR
		output wire        sram_LB_N,            //               .LB_N
		output wire        sram_UB_N,            //               .UB_N
		output wire        sram_CE_N,            //               .CE_N
		output wire        sram_OE_N,            //               .OE_N
		output wire        sram_WE_N,            //               .WE_N
		input  wire [17:0] switches_export,      //       switches.export
		output wire        vga_controller_CLK,   // vga_controller.CLK
		output wire        vga_controller_HS,    //               .HS
		output wire        vga_controller_VS,    //               .VS
		output wire        vga_controller_BLANK, //               .BLANK
		output wire        vga_controller_SYNC,  //               .SYNC
		output wire [7:0]  vga_controller_R,     //               .R
		output wire [7:0]  vga_controller_G,     //               .G
		output wire [7:0]  vga_controller_B      //               .B
	);

	wire         video_fifo_avalon_dc_buffer_source_valid;                           // video_fifo:stream_out_valid -> vga_controller:valid
	wire  [29:0] video_fifo_avalon_dc_buffer_source_data;                            // video_fifo:stream_out_data -> vga_controller:data
	wire         video_fifo_avalon_dc_buffer_source_ready;                           // vga_controller:ready -> video_fifo:stream_out_ready
	wire         video_fifo_avalon_dc_buffer_source_startofpacket;                   // video_fifo:stream_out_startofpacket -> vga_controller:startofpacket
	wire         video_fifo_avalon_dc_buffer_source_endofpacket;                     // video_fifo:stream_out_endofpacket -> vga_controller:endofpacket
	wire         pixel_buffer_dma_avalon_pixel_source_valid;                         // pixel_buffer_dma:stream_valid -> rgb_resampler:stream_in_valid
	wire  [15:0] pixel_buffer_dma_avalon_pixel_source_data;                          // pixel_buffer_dma:stream_data -> rgb_resampler:stream_in_data
	wire         pixel_buffer_dma_avalon_pixel_source_ready;                         // rgb_resampler:stream_in_ready -> pixel_buffer_dma:stream_ready
	wire         pixel_buffer_dma_avalon_pixel_source_startofpacket;                 // pixel_buffer_dma:stream_startofpacket -> rgb_resampler:stream_in_startofpacket
	wire         pixel_buffer_dma_avalon_pixel_source_endofpacket;                   // pixel_buffer_dma:stream_endofpacket -> rgb_resampler:stream_in_endofpacket
	wire         rgb_resampler_avalon_rgb_source_valid;                              // rgb_resampler:stream_out_valid -> scaler:stream_in_valid
	wire  [29:0] rgb_resampler_avalon_rgb_source_data;                               // rgb_resampler:stream_out_data -> scaler:stream_in_data
	wire         rgb_resampler_avalon_rgb_source_ready;                              // scaler:stream_in_ready -> rgb_resampler:stream_out_ready
	wire         rgb_resampler_avalon_rgb_source_startofpacket;                      // rgb_resampler:stream_out_startofpacket -> scaler:stream_in_startofpacket
	wire         rgb_resampler_avalon_rgb_source_endofpacket;                        // rgb_resampler:stream_out_endofpacket -> scaler:stream_in_endofpacket
	wire         scaler_avalon_scaler_source_valid;                                  // scaler:stream_out_valid -> video_fifo:stream_in_valid
	wire  [29:0] scaler_avalon_scaler_source_data;                                   // scaler:stream_out_data -> video_fifo:stream_in_data
	wire         scaler_avalon_scaler_source_ready;                                  // video_fifo:stream_in_ready -> scaler:stream_out_ready
	wire         scaler_avalon_scaler_source_startofpacket;                          // scaler:stream_out_startofpacket -> video_fifo:stream_in_startofpacket
	wire         scaler_avalon_scaler_source_endofpacket;                            // scaler:stream_out_endofpacket -> video_fifo:stream_in_endofpacket
	wire         sys_sdram_pll_0_sys_clk_clk;                                        // sys_sdram_pll_0:sys_clk_clk -> [address:clk, buttons:clk, din:clk, irq_mapper:clk, irq_synchronizer:sender_clk, jtag_uart:clk, leds:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, nios2_qsys_0:clk, onchip_memory:clk, pixel_buffer:clk, pixel_buffer_dma:clk, rgb_resampler:clk, rst_controller:clk, rst_controller_001:clk, scaler:clk, sdram:clk, switches:clk, video_fifo:clk_stream_in]
	wire         video_pll_0_vga_clk_clk;                                            // video_pll_0:vga_clk_clk -> [rst_controller_004:clk, vga_controller:clk, video_fifo:clk_stream_out]
	wire         pixel_buffer_dma_avalon_pixel_dma_master_waitrequest;               // mm_interconnect_0:pixel_buffer_dma_avalon_pixel_dma_master_waitrequest -> pixel_buffer_dma:master_waitrequest
	wire  [15:0] pixel_buffer_dma_avalon_pixel_dma_master_readdata;                  // mm_interconnect_0:pixel_buffer_dma_avalon_pixel_dma_master_readdata -> pixel_buffer_dma:master_readdata
	wire  [31:0] pixel_buffer_dma_avalon_pixel_dma_master_address;                   // pixel_buffer_dma:master_address -> mm_interconnect_0:pixel_buffer_dma_avalon_pixel_dma_master_address
	wire         pixel_buffer_dma_avalon_pixel_dma_master_read;                      // pixel_buffer_dma:master_read -> mm_interconnect_0:pixel_buffer_dma_avalon_pixel_dma_master_read
	wire         pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid;             // mm_interconnect_0:pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid -> pixel_buffer_dma:master_readdatavalid
	wire         pixel_buffer_dma_avalon_pixel_dma_master_lock;                      // pixel_buffer_dma:master_arbiterlock -> mm_interconnect_0:pixel_buffer_dma_avalon_pixel_dma_master_lock
	wire  [31:0] nios2_qsys_0_data_master_readdata;                                  // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                               // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                               // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [28:0] nios2_qsys_0_data_master_address;                                   // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                      // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_readdatavalid;                             // mm_interconnect_0:nios2_qsys_0_data_master_readdatavalid -> nios2_qsys_0:d_readdatavalid
	wire         nios2_qsys_0_data_master_write;                                     // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                 // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                           // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                        // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [28:0] nios2_qsys_0_instruction_master_address;                            // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                               // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         nios2_qsys_0_instruction_master_readdatavalid;                      // mm_interconnect_0:nios2_qsys_0_instruction_master_readdatavalid -> nios2_qsys_0:i_readdatavalid
	wire  [15:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdata;          // pixel_buffer:readdata -> mm_interconnect_0:pixel_buffer_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_address;           // mm_interconnect_0:pixel_buffer_avalon_sram_slave_address -> pixel_buffer:address
	wire         mm_interconnect_0_pixel_buffer_avalon_sram_slave_read;              // mm_interconnect_0:pixel_buffer_avalon_sram_slave_read -> pixel_buffer:read
	wire   [1:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_byteenable;        // mm_interconnect_0:pixel_buffer_avalon_sram_slave_byteenable -> pixel_buffer:byteenable
	wire         mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdatavalid;     // pixel_buffer:readdatavalid -> mm_interconnect_0:pixel_buffer_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_pixel_buffer_avalon_sram_slave_write;             // mm_interconnect_0:pixel_buffer_avalon_sram_slave_write -> pixel_buffer:write
	wire  [15:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_writedata;         // mm_interconnect_0:pixel_buffer_avalon_sram_slave_writedata -> pixel_buffer:writedata
	wire  [31:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata;   // pixel_buffer_dma:slave_readdata -> mm_interconnect_0:pixel_buffer_dma_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address;    // mm_interconnect_0:pixel_buffer_dma_avalon_control_slave_address -> pixel_buffer_dma:slave_address
	wire         mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read;       // mm_interconnect_0:pixel_buffer_dma_avalon_control_slave_read -> pixel_buffer_dma:slave_read
	wire   [3:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable; // mm_interconnect_0:pixel_buffer_dma_avalon_control_slave_byteenable -> pixel_buffer_dma:slave_byteenable
	wire         mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write;      // mm_interconnect_0:pixel_buffer_dma_avalon_control_slave_write -> pixel_buffer_dma:slave_write
	wire  [31:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata;  // mm_interconnect_0:pixel_buffer_dma_avalon_control_slave_writedata -> pixel_buffer_dma:slave_writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;             // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;          // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                 // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_buttons_avalon_parallel_port_slave_chipselect;    // mm_interconnect_0:buttons_avalon_parallel_port_slave_chipselect -> buttons:chipselect
	wire  [31:0] mm_interconnect_0_buttons_avalon_parallel_port_slave_readdata;      // buttons:readdata -> mm_interconnect_0:buttons_avalon_parallel_port_slave_readdata
	wire   [1:0] mm_interconnect_0_buttons_avalon_parallel_port_slave_address;       // mm_interconnect_0:buttons_avalon_parallel_port_slave_address -> buttons:address
	wire         mm_interconnect_0_buttons_avalon_parallel_port_slave_read;          // mm_interconnect_0:buttons_avalon_parallel_port_slave_read -> buttons:read
	wire   [3:0] mm_interconnect_0_buttons_avalon_parallel_port_slave_byteenable;    // mm_interconnect_0:buttons_avalon_parallel_port_slave_byteenable -> buttons:byteenable
	wire         mm_interconnect_0_buttons_avalon_parallel_port_slave_write;         // mm_interconnect_0:buttons_avalon_parallel_port_slave_write -> buttons:write
	wire  [31:0] mm_interconnect_0_buttons_avalon_parallel_port_slave_writedata;     // mm_interconnect_0:buttons_avalon_parallel_port_slave_writedata -> buttons:writedata
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;          // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest;       // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;           // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;              // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;             // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;         // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                      // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                        // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory_s1_address;                         // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                      // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                           // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                       // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                           // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                             // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                              // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_leds_s1_chipselect;                               // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                 // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                  // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                                    // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                              // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                                // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                             // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                 // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                    // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                              // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                           // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                   // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                               // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timer_0_s1_chipselect;                            // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                              // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                               // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                 // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                             // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire  [31:0] mm_interconnect_0_din_s1_readdata;                                  // din:readdata -> mm_interconnect_0:din_s1_readdata
	wire   [1:0] mm_interconnect_0_din_s1_address;                                   // mm_interconnect_0:din_s1_address -> din:address
	wire         mm_interconnect_0_address_s1_chipselect;                            // mm_interconnect_0:address_s1_chipselect -> address:chipselect
	wire  [31:0] mm_interconnect_0_address_s1_readdata;                              // address:readdata -> mm_interconnect_0:address_s1_readdata
	wire   [1:0] mm_interconnect_0_address_s1_address;                               // mm_interconnect_0:address_s1_address -> address:address
	wire         mm_interconnect_0_address_s1_write;                                 // mm_interconnect_0:address_s1_write -> address:write_n
	wire  [31:0] mm_interconnect_0_address_s1_writedata;                             // mm_interconnect_0:address_s1_writedata -> address:writedata
	wire         irq_mapper_receiver1_irq;                                           // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                             // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         irq_mapper_receiver0_irq;                                           // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                      // timer_0:irq -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [address:reset_n, din:reset_n, mm_interconnect_0:din_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> [buttons:reset, irq_mapper:reset, irq_synchronizer:sender_reset, jtag_uart:rst_n, leds:reset_n, mm_interconnect_0:pixel_buffer_dma_reset_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, onchip_memory:reset, pixel_buffer:reset, pixel_buffer_dma:reset, rgb_resampler:reset, rst_translator:in_reset, scaler:reset, sdram:reset_n, switches:reset_n, video_fifo:reset_stream_in]
	wire         rst_controller_001_reset_out_reset_req;                             // rst_controller_001:reset_req -> [nios2_qsys_0:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                         // nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_004:reset_in1]
	wire         rst_controller_002_reset_out_reset;                                 // rst_controller_002:reset_out -> [sys_sdram_pll_0:ref_reset_reset, video_pll_0:ref_reset_reset]
	wire         rst_controller_003_reset_out_reset;                                 // rst_controller_003:reset_out -> [irq_synchronizer:receiver_reset, mm_interconnect_0:timer_0_reset_reset_bridge_in_reset_reset, timer_0:reset_n]
	wire         rst_controller_004_reset_out_reset;                                 // rst_controller_004:reset_out -> [vga_controller:reset, video_fifo:reset_stream_out]

	nios_system_address address (
		.clk        (sys_sdram_pll_0_sys_clk_clk),             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_address_s1_readdata),   //                    .readdata
		.out_port   (address_export)                           // external_connection.export
	);

	nios_system_buttons buttons (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                                     //                        clk.clk
		.reset      (rst_controller_001_reset_out_reset),                              //                      reset.reset
		.address    (mm_interconnect_0_buttons_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_buttons_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_buttons_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_buttons_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_buttons_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_buttons_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_buttons_avalon_parallel_port_slave_readdata),   //                           .readdata
		.KEY        (buttons_export)                                                   //         external_interface.export
	);

	nios_system_din din (
		.clk      (sys_sdram_pll_0_sys_clk_clk),       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_din_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_din_s1_readdata), //                    .readdata
		.in_port  (din_export)                         // external_connection.export
	);

	nios_system_jtag_uart jtag_uart (
		.clk            (sys_sdram_pll_0_sys_clk_clk),                               //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	nios_system_leds leds (
		.clk        (sys_sdram_pll_0_sys_clk_clk),          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	nios_system_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (sys_sdram_pll_0_sys_clk_clk),                                  //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                          //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),                       //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_qsys_0_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_0_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	nios_system_onchip_memory onchip_memory (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                   //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)         //       .reset_req
	);

	nios_system_pixel_buffer pixel_buffer (
		.clk           (sys_sdram_pll_0_sys_clk_clk),                                    //                clk.clk
		.reset         (rst_controller_001_reset_out_reset),                             //              reset.reset
		.SRAM_DQ       (sram_DQ),                                                        // external_interface.export
		.SRAM_ADDR     (sram_ADDR),                                                      //                   .export
		.SRAM_LB_N     (sram_LB_N),                                                      //                   .export
		.SRAM_UB_N     (sram_UB_N),                                                      //                   .export
		.SRAM_CE_N     (sram_CE_N),                                                      //                   .export
		.SRAM_OE_N     (sram_OE_N),                                                      //                   .export
		.SRAM_WE_N     (sram_WE_N),                                                      //                   .export
		.address       (mm_interconnect_0_pixel_buffer_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_pixel_buffer_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_pixel_buffer_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_pixel_buffer_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_pixel_buffer_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	nios_system_pixel_buffer_dma pixel_buffer_dma (
		.clk                  (sys_sdram_pll_0_sys_clk_clk),                                        //                     clk.clk
		.reset                (rst_controller_001_reset_out_reset),                                 //                   reset.reset
		.master_readdatavalid (pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (pixel_buffer_dma_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (pixel_buffer_dma_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (pixel_buffer_dma_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (pixel_buffer_dma_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (pixel_buffer_dma_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_buffer_dma_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (pixel_buffer_dma_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (pixel_buffer_dma_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (pixel_buffer_dma_avalon_pixel_source_data)                           //                        .data
	);

	nios_system_rgb_resampler rgb_resampler (
		.clk                      (sys_sdram_pll_0_sys_clk_clk),                        //               clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                 //             reset.reset
		.stream_in_startofpacket  (pixel_buffer_dma_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixel_buffer_dma_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (pixel_buffer_dma_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (pixel_buffer_dma_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (pixel_buffer_dma_avalon_pixel_source_data),          //                  .data
		.stream_out_ready         (rgb_resampler_avalon_rgb_source_ready),              // avalon_rgb_source.ready
		.stream_out_startofpacket (rgb_resampler_avalon_rgb_source_startofpacket),      //                  .startofpacket
		.stream_out_endofpacket   (rgb_resampler_avalon_rgb_source_endofpacket),        //                  .endofpacket
		.stream_out_valid         (rgb_resampler_avalon_rgb_source_valid),              //                  .valid
		.stream_out_data          (rgb_resampler_avalon_rgb_source_data)                //                  .data
	);

	nios_system_scaler scaler (
		.clk                      (sys_sdram_pll_0_sys_clk_clk),                   //                  clk.clk
		.reset                    (rst_controller_001_reset_out_reset),            //                reset.reset
		.stream_in_startofpacket  (rgb_resampler_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (rgb_resampler_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (rgb_resampler_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (rgb_resampler_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (rgb_resampler_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (scaler_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (scaler_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (scaler_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (scaler_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (scaler_avalon_scaler_source_data)               //                     .data
	);

	nios_system_sdram sdram (
		.clk            (sys_sdram_pll_0_sys_clk_clk),              //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	nios_system_switches switches (
		.clk      (sys_sdram_pll_0_sys_clk_clk),            //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	nios_system_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_002_reset_out_reset), //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_0_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                      //    sdram_clk.clk
		.reset_source_reset ()                                    // reset_source.reset
	);

	nios_system_timer_0 timer_0 (
		.clk        (gameboy_clk_clk),                         //   clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)            //   irq.irq
	);

	nios_system_vga_controller vga_controller (
		.clk           (video_pll_0_vga_clk_clk),                          //                clk.clk
		.reset         (rst_controller_004_reset_out_reset),               //              reset.reset
		.data          (video_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_controller_CLK),                               // external_interface.export
		.VGA_HS        (vga_controller_HS),                                //                   .export
		.VGA_VS        (vga_controller_VS),                                //                   .export
		.VGA_BLANK     (vga_controller_BLANK),                             //                   .export
		.VGA_SYNC      (vga_controller_SYNC),                              //                   .export
		.VGA_R         (vga_controller_R),                                 //                   .export
		.VGA_G         (vga_controller_G),                                 //                   .export
		.VGA_B         (vga_controller_B)                                  //                   .export
	);

	nios_system_video_fifo video_fifo (
		.clk_stream_in            (sys_sdram_pll_0_sys_clk_clk),                      //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_001_reset_out_reset),               //         reset_stream_in.reset
		.clk_stream_out           (video_pll_0_vga_clk_clk),                          //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_004_reset_out_reset),               //        reset_stream_out.reset
		.stream_in_ready          (scaler_avalon_scaler_source_ready),                //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (scaler_avalon_scaler_source_startofpacket),        //                        .startofpacket
		.stream_in_endofpacket    (scaler_avalon_scaler_source_endofpacket),          //                        .endofpacket
		.stream_in_valid          (scaler_avalon_scaler_source_valid),                //                        .valid
		.stream_in_data           (scaler_avalon_scaler_source_data),                 //                        .data
		.stream_out_ready         (video_fifo_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_fifo_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (video_fifo_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (video_fifo_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (video_fifo_avalon_dc_buffer_source_data)           //                        .data
	);

	nios_system_video_pll_0 video_pll_0 (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_002_reset_out_reset), //    ref_reset.reset
		.vga_clk_clk        (video_pll_0_vga_clk_clk),            //      vga_clk.clk
		.reset_source_reset ()                                    // reset_source.reset
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.gameboy_clk_clk_clk                                    (gameboy_clk_clk),                                                    //                              gameboy_clk_clk.clk
		.sys_sdram_pll_0_sys_clk_clk                            (sys_sdram_pll_0_sys_clk_clk),                                        //                      sys_sdram_pll_0_sys_clk.clk
		.din_reset_reset_bridge_in_reset_reset                  (rst_controller_reset_out_reset),                                     //              din_reset_reset_bridge_in_reset.reset
		.pixel_buffer_dma_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                                 // pixel_buffer_dma_reset_reset_bridge_in_reset.reset
		.timer_0_reset_reset_bridge_in_reset_reset              (rst_controller_003_reset_out_reset),                                 //          timer_0_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                       (nios2_qsys_0_data_master_address),                                   //                     nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest                   (nios2_qsys_0_data_master_waitrequest),                               //                                             .waitrequest
		.nios2_qsys_0_data_master_byteenable                    (nios2_qsys_0_data_master_byteenable),                                //                                             .byteenable
		.nios2_qsys_0_data_master_read                          (nios2_qsys_0_data_master_read),                                      //                                             .read
		.nios2_qsys_0_data_master_readdata                      (nios2_qsys_0_data_master_readdata),                                  //                                             .readdata
		.nios2_qsys_0_data_master_readdatavalid                 (nios2_qsys_0_data_master_readdatavalid),                             //                                             .readdatavalid
		.nios2_qsys_0_data_master_write                         (nios2_qsys_0_data_master_write),                                     //                                             .write
		.nios2_qsys_0_data_master_writedata                     (nios2_qsys_0_data_master_writedata),                                 //                                             .writedata
		.nios2_qsys_0_data_master_debugaccess                   (nios2_qsys_0_data_master_debugaccess),                               //                                             .debugaccess
		.nios2_qsys_0_instruction_master_address                (nios2_qsys_0_instruction_master_address),                            //              nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest            (nios2_qsys_0_instruction_master_waitrequest),                        //                                             .waitrequest
		.nios2_qsys_0_instruction_master_read                   (nios2_qsys_0_instruction_master_read),                               //                                             .read
		.nios2_qsys_0_instruction_master_readdata               (nios2_qsys_0_instruction_master_readdata),                           //                                             .readdata
		.nios2_qsys_0_instruction_master_readdatavalid          (nios2_qsys_0_instruction_master_readdatavalid),                      //                                             .readdatavalid
		.pixel_buffer_dma_avalon_pixel_dma_master_address       (pixel_buffer_dma_avalon_pixel_dma_master_address),                   //     pixel_buffer_dma_avalon_pixel_dma_master.address
		.pixel_buffer_dma_avalon_pixel_dma_master_waitrequest   (pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),               //                                             .waitrequest
		.pixel_buffer_dma_avalon_pixel_dma_master_read          (pixel_buffer_dma_avalon_pixel_dma_master_read),                      //                                             .read
		.pixel_buffer_dma_avalon_pixel_dma_master_readdata      (pixel_buffer_dma_avalon_pixel_dma_master_readdata),                  //                                             .readdata
		.pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid (pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),             //                                             .readdatavalid
		.pixel_buffer_dma_avalon_pixel_dma_master_lock          (pixel_buffer_dma_avalon_pixel_dma_master_lock),                      //                                             .lock
		.address_s1_address                                     (mm_interconnect_0_address_s1_address),                               //                                   address_s1.address
		.address_s1_write                                       (mm_interconnect_0_address_s1_write),                                 //                                             .write
		.address_s1_readdata                                    (mm_interconnect_0_address_s1_readdata),                              //                                             .readdata
		.address_s1_writedata                                   (mm_interconnect_0_address_s1_writedata),                             //                                             .writedata
		.address_s1_chipselect                                  (mm_interconnect_0_address_s1_chipselect),                            //                                             .chipselect
		.buttons_avalon_parallel_port_slave_address             (mm_interconnect_0_buttons_avalon_parallel_port_slave_address),       //           buttons_avalon_parallel_port_slave.address
		.buttons_avalon_parallel_port_slave_write               (mm_interconnect_0_buttons_avalon_parallel_port_slave_write),         //                                             .write
		.buttons_avalon_parallel_port_slave_read                (mm_interconnect_0_buttons_avalon_parallel_port_slave_read),          //                                             .read
		.buttons_avalon_parallel_port_slave_readdata            (mm_interconnect_0_buttons_avalon_parallel_port_slave_readdata),      //                                             .readdata
		.buttons_avalon_parallel_port_slave_writedata           (mm_interconnect_0_buttons_avalon_parallel_port_slave_writedata),     //                                             .writedata
		.buttons_avalon_parallel_port_slave_byteenable          (mm_interconnect_0_buttons_avalon_parallel_port_slave_byteenable),    //                                             .byteenable
		.buttons_avalon_parallel_port_slave_chipselect          (mm_interconnect_0_buttons_avalon_parallel_port_slave_chipselect),    //                                             .chipselect
		.din_s1_address                                         (mm_interconnect_0_din_s1_address),                                   //                                       din_s1.address
		.din_s1_readdata                                        (mm_interconnect_0_din_s1_readdata),                                  //                                             .readdata
		.jtag_uart_avalon_jtag_slave_address                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),              //                  jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                //                                             .write
		.jtag_uart_avalon_jtag_slave_read                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                 //                                             .read
		.jtag_uart_avalon_jtag_slave_readdata                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),             //                                             .readdata
		.jtag_uart_avalon_jtag_slave_writedata                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),            //                                             .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),          //                                             .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),           //                                             .chipselect
		.leds_s1_address                                        (mm_interconnect_0_leds_s1_address),                                  //                                      leds_s1.address
		.leds_s1_write                                          (mm_interconnect_0_leds_s1_write),                                    //                                             .write
		.leds_s1_readdata                                       (mm_interconnect_0_leds_s1_readdata),                                 //                                             .readdata
		.leds_s1_writedata                                      (mm_interconnect_0_leds_s1_writedata),                                //                                             .writedata
		.leds_s1_chipselect                                     (mm_interconnect_0_leds_s1_chipselect),                               //                                             .chipselect
		.nios2_qsys_0_jtag_debug_module_address                 (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),           //               nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write                   (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),             //                                             .write
		.nios2_qsys_0_jtag_debug_module_read                    (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),              //                                             .read
		.nios2_qsys_0_jtag_debug_module_readdata                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),          //                                             .readdata
		.nios2_qsys_0_jtag_debug_module_writedata               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),         //                                             .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),        //                                             .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest),       //                                             .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess),       //                                             .debugaccess
		.onchip_memory_s1_address                               (mm_interconnect_0_onchip_memory_s1_address),                         //                             onchip_memory_s1.address
		.onchip_memory_s1_write                                 (mm_interconnect_0_onchip_memory_s1_write),                           //                                             .write
		.onchip_memory_s1_readdata                              (mm_interconnect_0_onchip_memory_s1_readdata),                        //                                             .readdata
		.onchip_memory_s1_writedata                             (mm_interconnect_0_onchip_memory_s1_writedata),                       //                                             .writedata
		.onchip_memory_s1_byteenable                            (mm_interconnect_0_onchip_memory_s1_byteenable),                      //                                             .byteenable
		.onchip_memory_s1_chipselect                            (mm_interconnect_0_onchip_memory_s1_chipselect),                      //                                             .chipselect
		.onchip_memory_s1_clken                                 (mm_interconnect_0_onchip_memory_s1_clken),                           //                                             .clken
		.pixel_buffer_avalon_sram_slave_address                 (mm_interconnect_0_pixel_buffer_avalon_sram_slave_address),           //               pixel_buffer_avalon_sram_slave.address
		.pixel_buffer_avalon_sram_slave_write                   (mm_interconnect_0_pixel_buffer_avalon_sram_slave_write),             //                                             .write
		.pixel_buffer_avalon_sram_slave_read                    (mm_interconnect_0_pixel_buffer_avalon_sram_slave_read),              //                                             .read
		.pixel_buffer_avalon_sram_slave_readdata                (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdata),          //                                             .readdata
		.pixel_buffer_avalon_sram_slave_writedata               (mm_interconnect_0_pixel_buffer_avalon_sram_slave_writedata),         //                                             .writedata
		.pixel_buffer_avalon_sram_slave_byteenable              (mm_interconnect_0_pixel_buffer_avalon_sram_slave_byteenable),        //                                             .byteenable
		.pixel_buffer_avalon_sram_slave_readdatavalid           (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdatavalid),     //                                             .readdatavalid
		.pixel_buffer_dma_avalon_control_slave_address          (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address),    //        pixel_buffer_dma_avalon_control_slave.address
		.pixel_buffer_dma_avalon_control_slave_write            (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write),      //                                             .write
		.pixel_buffer_dma_avalon_control_slave_read             (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read),       //                                             .read
		.pixel_buffer_dma_avalon_control_slave_readdata         (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata),   //                                             .readdata
		.pixel_buffer_dma_avalon_control_slave_writedata        (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata),  //                                             .writedata
		.pixel_buffer_dma_avalon_control_slave_byteenable       (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable), //                                             .byteenable
		.sdram_s1_address                                       (mm_interconnect_0_sdram_s1_address),                                 //                                     sdram_s1.address
		.sdram_s1_write                                         (mm_interconnect_0_sdram_s1_write),                                   //                                             .write
		.sdram_s1_read                                          (mm_interconnect_0_sdram_s1_read),                                    //                                             .read
		.sdram_s1_readdata                                      (mm_interconnect_0_sdram_s1_readdata),                                //                                             .readdata
		.sdram_s1_writedata                                     (mm_interconnect_0_sdram_s1_writedata),                               //                                             .writedata
		.sdram_s1_byteenable                                    (mm_interconnect_0_sdram_s1_byteenable),                              //                                             .byteenable
		.sdram_s1_readdatavalid                                 (mm_interconnect_0_sdram_s1_readdatavalid),                           //                                             .readdatavalid
		.sdram_s1_waitrequest                                   (mm_interconnect_0_sdram_s1_waitrequest),                             //                                             .waitrequest
		.sdram_s1_chipselect                                    (mm_interconnect_0_sdram_s1_chipselect),                              //                                             .chipselect
		.switches_s1_address                                    (mm_interconnect_0_switches_s1_address),                              //                                  switches_s1.address
		.switches_s1_readdata                                   (mm_interconnect_0_switches_s1_readdata),                             //                                             .readdata
		.timer_0_s1_address                                     (mm_interconnect_0_timer_0_s1_address),                               //                                   timer_0_s1.address
		.timer_0_s1_write                                       (mm_interconnect_0_timer_0_s1_write),                                 //                                             .write
		.timer_0_s1_readdata                                    (mm_interconnect_0_timer_0_s1_readdata),                              //                                             .readdata
		.timer_0_s1_writedata                                   (mm_interconnect_0_timer_0_s1_writedata),                             //                                             .writedata
		.timer_0_s1_chipselect                                  (mm_interconnect_0_timer_0_s1_chipselect)                             //                                             .chipselect
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (sys_sdram_pll_0_sys_clk_clk),        //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)              //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (gameboy_clk_clk),                    //       receiver_clk.clk
		.sender_clk     (sys_sdram_pll_0_sys_clk_clk),        //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (gameboy_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (video_pll_0_vga_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
